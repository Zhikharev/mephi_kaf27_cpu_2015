`include "cpu_interface.sv"
`include "model_pkg.sv"
`include "transaction.sv"
`include "topmodule.sv"
`include "inst_driver.sv"
`include "inst_monitor.sv"
`include "data_monitor.sv"
`include "data_driver.sv"
`include "environment.sv"
//`include "testcase.sv"
