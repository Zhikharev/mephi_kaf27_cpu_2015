`ifndef TRANZACTION
`define TRANZACTION


class tranz 
        rand 














`endif 
