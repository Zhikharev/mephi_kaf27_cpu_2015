/*
`include "cpu_interface.sv"
`include "model_pkg.sv"
`include "transaction.sv"
`include "inst_driver.sv"
`include "inst_monitor.sv"
`include "data_monitor.sv"
`include "data_driver.sv"
`include "environment.sv"
`include "testcase.sv"
`include "topmodule.sv" 
*/
`include "my_cpu_interface.sv"
//`include "my_transaction.sv"
`include "my_3transaction.sv"
`include "my_instr_driver.sv"
`include "ideal_cpu.sv"
`include "my_scorebord.sv"
`include "my_mem.sv"
`include "my_environment.sv"
`include "my_testcase.sv"
`include "my_topmodule.sv"
