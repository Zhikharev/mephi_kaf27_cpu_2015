package model;

	import "DPI-C" function void test_sv_c_communication(input int val);
	import "DPI-C" function  decode(int,int);//int instr, int verbosity
	import "DPI-C" function init_memory();
    import "DPI-C" function set_memory(int,int);//addr data
    import "DPI-C" function get_memory(int); //addr 
    import "DPI-C" function ADD(int,int,int);//rs rt rd
    import "DPI-C" function ADDI(int,int,int);
    import "DPI-C" function OR(int,int,int);
    import "DPI-C" function AND(int,int,int);
    import "DPI-C" function XOR(int,int,int);
    import "DPI-C" function NOR(int,int,int);
    import "DPI-C" function SLL(int,int,int);
    import "DPI-C" function ROT(int,int,int);
    import "DPI-C" function BNE(int,int,int);
    import "DPI-C" function LDL(int);
    import "DPI-C" function LDH(int);
    import "DPI-C" function STL(int);
    import "DPI-C" function STH(int);
    import "DPI-C" function JMP(int);
    import "DPI-C" function JAL(int);
    import "DPI-C" function JR(int);
    import "DPI-C" function JARL(int);
    import "DPI-C" function NOP();
    import "DPI-C" function aiireg(int); //int verbosity
    import "DPI-C" function statistic(int); //int verbosity 
    import "DPI-C" function write_resalt();
 

    
    
endpackage
