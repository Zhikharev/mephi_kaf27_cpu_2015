`include "defines.v"
`include "chu_dpi.sv"
`include "chu_pad_interface.sv"
`include "chu_pad_packet.sv"
`include "chu_pad_driver.sv"
`include "chu_pad_monitor.sv" 
`include "chu_pad_scoreboard.sv"
`include "chu_pad_environment.sv"
`include "chu_pad_testcase.sv"
`include "chu_pad_top.sv"
