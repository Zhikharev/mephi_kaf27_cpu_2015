`ifndef TESTCASE
`define TESCASE
//$display("testcase was read");













`endif
