`include "cpu_interface.sv"
//`include "model_pkg.sv"
`include "transaction.sv"
`include "topmodule.sv"
`include "driver.sv"
