
import "DPI-C" function void md5_align(output bit [31:0] ext[64], input string mes, input int size_from_sv);
import "DPI-C" function  void sha1_align(output bit [31:0] ext[64], input string mes);
