`ifndef MONITOR
`define MONITOR
class monitor;
    virtual wishbone mon_int;
    virtual control mon_control;
    //mailbox #()




















`endif
