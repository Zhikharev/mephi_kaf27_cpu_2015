package model;

	import "DPI-C" function void test_sv_c_communication(input int val);

endpackage