`ifndef DATA_MONITOR
`define DATA_MONITOR

class data_monitor




endclass








`endif
