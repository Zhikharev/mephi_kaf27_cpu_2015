`include "cpu_interface.sv"
`include "transaction.sv"
`include "topmodule.sv"
