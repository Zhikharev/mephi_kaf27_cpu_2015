`ifdef ENVIRONMENT
`define ENVIRONMENT


class environment
        virtual cpu_int vir_cpu_int;
        
        function new 













`endif
