module cpu (
	input CLK_I,
	input RTS_I,
	input[15:0] ADR_I,
	input [15:0] DAT_I,
	output[15:0] ADR_O,
	output [15:0] DAT_O
	);
endmodule
