`include "cpu_interface.sv"
`include "model_pkg.sv"
`include "transaction.sv"
`include "topmodule.sv"
//`include "driver.sv"
`include "monitor.sv"
`include "environment.sv"
