`include "cpu_interface.sv"
`include "topmodule.sv"